library ieee;
use ieee.std_logic_1164.all;

entity mux is
end mux;

architecture behavioral of mux is

begin

end architecture;